package mips_pkg;
    parameter PC_WIDTH       = 32;
    parameter INSTR_WITDTH   = 32;
    parameter DATA_MEM_WIDTH = 32;
    parameter ALU_CTRL_WIDTH = 3; 
endpackage