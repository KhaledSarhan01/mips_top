////////////////////////////////////////////////
///// Project   : mips_top             
///// Created on: 2025-11-20                   
////////////////////////////////////////////////

module mips_top (
// Clock and active low Asynchronous Reset
    input logic clk,rst_n 
// Signals    
    
);
// Enter your code here
// THIS IS DUMMY CODE
    
endmodule
